module nand_gate(Y,A,B);
	input A,B;
	output Y;
	nand (Y,A,B);
endmodule
